// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
// Created on Sun Feb 25 15:57:28 2018

// synthesis message_off 10175

`timescale 1ns/1ns

module SquareWaveGenerator (
    clock,reset,a,b,
    out1);

    input clock;
    input reset;
    input a;
    input b;
    tri0 reset;
    tri0 a;
    tri0 b;
    output out1;
    reg out1;
    reg reg_out1;
    reg [1:0] fstate;
    reg [1:0] reg_fstate;
    parameter state1=0,state2=1;

    initial
    begin
        reg_out1 <= 1'b0;
    end

    always @(posedge clock or posedge reset)
    begin
        if (reset) begin
            fstate <= state1;
        end
        else begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or a or b or reg_out1)
    begin
        reg_out1 <= 1'b0;
        out1 <= 1'b0;
        case (fstate)
            state1: begin
                if (a)
                    reg_fstate <= state2;
                // Inserting 'else' block to prevent latch inference
                else
                    reg_fstate <= state1;

                reg_out1 <= (a | b);
            end
            state2: begin
                if (~(a))
                    reg_fstate <= state1;
                // Inserting 'else' block to prevent latch inference
                else
                    reg_fstate <= state2;

                reg_out1 <= a;
            end
            default: begin
                reg_out1 <= 1'bx;
                $display ("Reach undefined state");
            end
        endcase
        out1 <= reg_out1;
    end
endmodule // SquareWaveGenerator
